class fifo_model extends model #(fifo_packet);
    function packet_t_queue get_expected_packet(fifo_packet input_packet);
        fifo_packet             expected_values[$];
        expected_values[0]    = input_packet;
        return expected_values;
    endfunction
endclass: fifo_model